`ifndef HVSYNC
`define HVSYNC

/*
Video sync generator, used to drive a simulated CRT.
To use:
- Wire the hsync and vsync signals to top level outputs
- Add a 3-bit (or more) "rgb" output to the top level
*/

module hvsync_generator(clk, reset, hsync, vsync, display_on, hpos, vpos);

  input clk;
  input reset;
  output reg hsync, vsync;
  output display_on;
  reg [8:0] hpos_internal;
  reg [8:0] vpos_internal;
  output [8:0] hpos;
  output [8:0] vpos;
  
  assign hpos = hpos_internal;
  assign vpos = vpos_internal;
  
  // sync RAM adjustment
  assign hpos = hpos_internal >= H_SYNC_START ? 0 : hpos_internal + 1;
  assign vpos = vpos_internal >= V_SYNC_START ? 0 :
    hpos_internal >= H_SYNC_START ? vpos_internal + 1 : vpos_internal;
  
  // declarations for TV-simulator sync parameters
  // horizontal constants
  parameter H_DISPLAY       = 256; // horizontal display width
  parameter H_BACK          =  23; // horizontal left border (back porch)
  parameter H_FRONT         =   7; // horizontal right border (front porch)
  parameter H_SYNC          =  23; // horizontal sync width
  // vertical constants
  parameter V_DISPLAY       = 240; // vertical display height
  parameter V_TOP           =   5; // vertical top border
  parameter V_BOTTOM        =  14; // vertical bottom border
  parameter V_SYNC          =   3; // vertical sync # lines
  // derived constants
  parameter H_SYNC_START    = H_DISPLAY + H_FRONT;
  parameter H_SYNC_END      = H_DISPLAY + H_FRONT + H_SYNC - 1;
  parameter H_MAX           = H_DISPLAY + H_BACK + H_FRONT + H_SYNC - 1;
  parameter V_SYNC_START    = V_DISPLAY + V_BOTTOM;
  parameter V_SYNC_END      = V_DISPLAY + V_BOTTOM + V_SYNC - 1;
  parameter V_MAX           = V_DISPLAY + V_TOP + V_BOTTOM + V_SYNC - 1;

  wire hmaxxed = (hpos_internal == H_MAX) || reset;    // set when hpos is maximum
  wire vmaxxed = (vpos_internal == V_MAX) || reset;    // set when vpos is maximum
  
  // horizontal position counter
  always @(posedge clk)
  begin
    hsync <= (hpos_internal>=H_SYNC_START && hpos_internal<=H_SYNC_END);
    if(hmaxxed)
      hpos_internal <= 0;
    else
      hpos_internal <= hpos_internal + 1;
  end

  // vertical position counter
  always @(posedge clk)
  begin
    vsync <= (vpos_internal>=V_SYNC_START && vpos_internal<=V_SYNC_END);
    if(hmaxxed)
      if (vmaxxed)
        vpos_internal <= 0;
      else
        vpos_internal <= vpos_internal + 1;
  end
  
  // display_on is set when beam is in "safe" visible frame
  assign display_on = (hpos_internal<H_DISPLAY) && (vpos_internal<V_DISPLAY);

endmodule

`endif
